module And_Gate(a,b,c);

input a,b;
output c;

assign c = a&b;

endmodule